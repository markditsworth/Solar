P. Basso: Switched-Mode Power Supplies, 2008, Chapter 1
* boost-converter
* Fig. 1-27

.control
set xtrtol=2
*save @V1[i] @V1[p] @Vin[i] @Vin[p] @Rload[i] @Rload[p]
*save @L1[i] @C1[i] @D1[id] @D1[p] @Resr[i] @Resr[p]
save 1 3 2 V(4) V(5) I(Vin)
run
plot v(1)
.endc

.TRAN 0.1u 1m 0 100n
.OPTIONS method=GEAR
.OPTIONS reltol=0.01
.PRINT  TRAN Vout

asw1 2 (0 3) switch3
.model switch3 aswitch(cntl_off=2.0 cntl_on=3.0 r_off=1e6
+ r_on=10m log=TRUE)

L1 4 3 1u
V1 2 0 PULSE 0 5 0 1n 1n 2.45u 8.33u 
Vin 4 0 DC=12
Rload 1 0 1
C1 1 5 3000u
D1 3 1 1n5818
.MODEL 1n5818 d AF=1 BV=30 CJO=1.98376e-10 EG=0.6 FC=0.5
+ IBV=0.001 IS=4.4214e-05 KF=0 M=0.54046 N=1.37435
+ RS=0.0531374 TT=2.6273e-08 VJ=1.5 XTI=0.5
Resr 5 0 100m
.END 
